`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:07:02 10/31/2020 
// Design Name: 
// Module Name:    HALF_ADDER_ 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module HALF_ADDER_(a,b,sum
    );
input a,b;
output sum;
xor(sum,a,b);
endmodule
